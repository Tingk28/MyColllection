module Vending(
    clk,
    rst,
    DI,
    MI,
    sel,
    re,
    MO,
    PO
);
    input clk;
    input rst;
    input [7:0] DI;
    input [7:0] MI;
    input [1:0] sel;
    input       re;
    output [7:0] MO;
    output [1:0] PO;

    // Complete this part by yourself

endmodule